`include "myfilter.svh"
import myfilter_pkg::*;

module dpc
  
  (input logic clk,
   input logic rst_n,
   input logic ul_in,
   input logic dl_in, 
   input logic extready_in, 
   output      dp_cmd_t cmd_out );

   
endmodule


