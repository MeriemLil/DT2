`include "myfilter.svh"
import myfilter_pkg::*;

module i2c_ctr
  
  (input logic clk,
   input logic 	rst_n,
   input logic 	clr_in,
   input logic 	next_in,
   input logic 	byteen_in, 
   output logic byteok_out,
   output logic frameok_out   
   );

   
endmodule


