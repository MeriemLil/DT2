`include "myfilter.svh"
import myfilter_pkg::*;

module reset_sync
  
  (input logic clk,
   input logic rst_n,
   output logic srst_n   
   );

   
endmodule

