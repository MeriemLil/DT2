`include "myfilter.svh"
import myfilter_pkg::*;

module i2c_srg
  
  (input logic clk,
   input logic 	     rst_n,
   input logic 	     clr_in,
   input logic 	     next_in,
   input logic 	     bit_in,
   output logic      bit_out,
   output logic      addrok_out
   );

  
endmodule


